* SPICE3 file created from XORinv.ext - technology: scmos

.include TSMC_180nm.txt

vdd vdd gnd 2.0V

.option scale=0.09u

Vin1 a gnd pulse(0 2.0 0 0.01p 0.01p 10n 20n)
Vin2 b gnd pulse(0 2.0 0 0.01p 0.01p 20n 40n)

M1000 out b vdd w_n25_63# CMOSP w=8 l=2
+  ad=40 pd=26 as=228 ps=138
M1001 out b gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=150 ps=64
M1002 NOT_1/out a vdd NOT_1/w_0_0# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1003 NOT_1/out a gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=20 ps=18
M1004 vdd b XOR_0/a_n5_3# XOR_0/w_n57_n3# CMOSP w=9 l=4
+  ad=0 pd=0 as=162 ps=54
M1005 gnd a XOR_0/a_n41_n54# gnd CMOSN w=13 l=4
+  ad=0 pd=0 as=468 ps=124
M1006 outout b XOR_0/a_n41_n54# gnd CMOSN w=13 l=4
+  ad=624 pd=148 as=0 ps=0
M1007 XOR_0/a_n41_n54# out outout gnd CMOSN w=13 l=4
+  ad=0 pd=0 as=0 ps=0
M1008 XOR_0/a_n41_n54# NOT_1/out gnd gnd CMOSN w=13 l=4
+  ad=0 pd=0 as=0 ps=0
M1009 XOR_0/a_n5_3# NOT_1/out outout XOR_0/w_n57_n3# CMOSP w=9 l=4
+  ad=0 pd=0 as=90 ps=38
M1010 XOR_0/a_n41_3# out vdd XOR_0/w_n57_n3# CMOSP w=9 l=4
+  ad=162 pd=54 as=0 ps=0
M1011 outout a XOR_0/a_n41_3# XOR_0/w_n57_n3# CMOSP w=9 l=4
+  ad=0 pd=0 as=0 ps=0

.control
tran 1n 160n
plot v(a)
plot v(b)
plot v(outout)
.endc
.end