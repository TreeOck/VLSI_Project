magic
tech scmos
timestamp 1638835252
<< nwell >>
rect 30 -105 54 -85
rect -5 -168 81 -147
rect -47 -188 -23 -168
rect -12 -289 50 -268
rect 59 -319 83 -299
rect 30 -388 54 -368
rect -5 -451 81 -430
rect -47 -471 -23 -451
rect -12 -572 50 -551
rect 59 -602 83 -582
rect 30 -660 54 -640
rect -5 -723 81 -702
rect -47 -743 -23 -723
rect -12 -844 50 -823
rect 59 -874 83 -854
<< ntransistor >>
rect 41 -117 43 -113
rect -36 -200 -34 -196
rect 7 -219 11 -206
rect 29 -219 33 -206
rect 43 -219 47 -206
rect 65 -219 69 -206
rect 7 -327 12 -318
rect 25 -327 30 -318
rect 70 -331 72 -327
rect 41 -400 43 -396
rect -36 -483 -34 -479
rect 7 -502 11 -489
rect 29 -502 33 -489
rect 43 -502 47 -489
rect 65 -502 69 -489
rect 7 -610 12 -601
rect 25 -610 30 -601
rect 70 -614 72 -610
rect 41 -672 43 -668
rect -36 -755 -34 -751
rect 7 -774 11 -761
rect 29 -774 33 -761
rect 43 -774 47 -761
rect 65 -774 69 -761
rect 7 -882 12 -873
rect 25 -882 30 -873
rect 70 -886 72 -882
<< ptransistor >>
rect 41 -99 43 -91
rect 7 -162 11 -153
rect 29 -162 33 -153
rect 43 -162 47 -153
rect 65 -162 69 -153
rect -36 -182 -34 -174
rect 7 -283 12 -274
rect 25 -283 30 -274
rect 70 -313 72 -305
rect 41 -382 43 -374
rect 7 -445 11 -436
rect 29 -445 33 -436
rect 43 -445 47 -436
rect 65 -445 69 -436
rect -36 -465 -34 -457
rect 7 -566 12 -557
rect 25 -566 30 -557
rect 70 -596 72 -588
rect 41 -654 43 -646
rect 7 -717 11 -708
rect 29 -717 33 -708
rect 43 -717 47 -708
rect 65 -717 69 -708
rect -36 -737 -34 -729
rect 7 -838 12 -829
rect 25 -838 30 -829
rect 70 -868 72 -860
<< ndiffusion >>
rect 40 -117 41 -113
rect 43 -117 44 -113
rect -37 -200 -36 -196
rect -34 -200 -33 -196
rect -15 -217 -8 -206
rect 0 -217 7 -206
rect -15 -219 7 -217
rect 11 -217 12 -206
rect 16 -208 29 -206
rect 16 -217 24 -208
rect 11 -219 24 -217
rect 28 -219 29 -208
rect 33 -210 43 -206
rect 33 -219 34 -210
rect 42 -219 43 -210
rect 47 -217 48 -206
rect 52 -208 65 -206
rect 52 -217 60 -208
rect 47 -219 60 -217
rect 64 -219 65 -208
rect 69 -217 80 -206
rect 88 -217 95 -206
rect 69 -219 95 -217
rect -3 -320 7 -318
rect -3 -327 -2 -320
rect 4 -327 7 -320
rect 12 -327 25 -318
rect 30 -325 33 -318
rect 38 -325 45 -318
rect 30 -327 45 -325
rect 69 -331 70 -327
rect 72 -331 73 -327
rect 40 -400 41 -396
rect 43 -400 44 -396
rect -37 -483 -36 -479
rect -34 -483 -33 -479
rect -15 -500 -8 -489
rect 0 -500 7 -489
rect -15 -502 7 -500
rect 11 -500 12 -489
rect 16 -491 29 -489
rect 16 -500 24 -491
rect 11 -502 24 -500
rect 28 -502 29 -491
rect 33 -493 43 -489
rect 33 -502 34 -493
rect 42 -502 43 -493
rect 47 -500 48 -489
rect 52 -491 65 -489
rect 52 -500 60 -491
rect 47 -502 60 -500
rect 64 -502 65 -491
rect 69 -500 80 -489
rect 88 -500 95 -489
rect 69 -502 95 -500
rect -3 -603 7 -601
rect -3 -610 -2 -603
rect 4 -610 7 -603
rect 12 -610 25 -601
rect 30 -608 33 -601
rect 38 -608 45 -601
rect 30 -610 45 -608
rect 69 -614 70 -610
rect 72 -614 73 -610
rect 40 -672 41 -668
rect 43 -672 44 -668
rect -37 -755 -36 -751
rect -34 -755 -33 -751
rect -15 -772 -8 -761
rect 0 -772 7 -761
rect -15 -774 7 -772
rect 11 -772 12 -761
rect 16 -763 29 -761
rect 16 -772 24 -763
rect 11 -774 24 -772
rect 28 -774 29 -763
rect 33 -765 43 -761
rect 33 -774 34 -765
rect 42 -774 43 -765
rect 47 -772 48 -761
rect 52 -763 65 -761
rect 52 -772 60 -763
rect 47 -774 60 -772
rect 64 -774 65 -763
rect 69 -772 80 -761
rect 88 -772 95 -761
rect 69 -774 95 -772
rect -3 -875 7 -873
rect -3 -882 -2 -875
rect 4 -882 7 -875
rect 12 -882 25 -873
rect 30 -880 33 -873
rect 38 -880 45 -873
rect 30 -882 45 -880
rect 69 -886 70 -882
rect 72 -886 73 -882
<< pdiffusion >>
rect 40 -99 41 -91
rect 43 -99 44 -91
rect 1 -159 2 -153
rect 6 -159 7 -153
rect 1 -162 7 -159
rect 11 -162 29 -153
rect 33 -154 43 -153
rect 33 -162 34 -154
rect 42 -162 43 -154
rect 47 -162 65 -153
rect 69 -159 70 -153
rect 74 -159 75 -153
rect 69 -162 75 -159
rect -37 -182 -36 -174
rect -34 -182 -33 -174
rect -5 -279 -2 -274
rect 3 -279 7 -274
rect -5 -283 7 -279
rect 12 -277 25 -274
rect 12 -283 16 -277
rect 22 -283 25 -277
rect 30 -279 36 -274
rect 41 -279 43 -274
rect 30 -283 43 -279
rect 69 -313 70 -305
rect 72 -313 73 -305
rect 40 -382 41 -374
rect 43 -382 44 -374
rect 1 -442 2 -436
rect 6 -442 7 -436
rect 1 -445 7 -442
rect 11 -445 29 -436
rect 33 -437 43 -436
rect 33 -445 34 -437
rect 42 -445 43 -437
rect 47 -445 65 -436
rect 69 -442 70 -436
rect 74 -442 75 -436
rect 69 -445 75 -442
rect -37 -465 -36 -457
rect -34 -465 -33 -457
rect -5 -562 -2 -557
rect 3 -562 7 -557
rect -5 -566 7 -562
rect 12 -560 25 -557
rect 12 -566 16 -560
rect 22 -566 25 -560
rect 30 -562 36 -557
rect 41 -562 43 -557
rect 30 -566 43 -562
rect 69 -596 70 -588
rect 72 -596 73 -588
rect 40 -654 41 -646
rect 43 -654 44 -646
rect 1 -714 2 -708
rect 6 -714 7 -708
rect 1 -717 7 -714
rect 11 -717 29 -708
rect 33 -709 43 -708
rect 33 -717 34 -709
rect 42 -717 43 -709
rect 47 -717 65 -708
rect 69 -714 70 -708
rect 74 -714 75 -708
rect 69 -717 75 -714
rect -37 -737 -36 -729
rect -34 -737 -33 -729
rect -5 -834 -2 -829
rect 3 -834 7 -829
rect -5 -838 7 -834
rect 12 -832 25 -829
rect 12 -838 16 -832
rect 22 -838 25 -832
rect 30 -834 36 -829
rect 41 -834 43 -829
rect 30 -838 43 -834
rect 69 -868 70 -860
rect 72 -868 73 -860
<< ndcontact >>
rect 36 -117 40 -113
rect 44 -117 48 -113
rect -41 -200 -37 -196
rect -33 -200 -29 -196
rect -8 -217 0 -206
rect 12 -217 16 -206
rect 24 -219 28 -208
rect 34 -219 42 -210
rect 48 -217 52 -206
rect 60 -219 64 -208
rect 80 -217 88 -206
rect -2 -327 4 -320
rect 33 -325 38 -318
rect 65 -331 69 -327
rect 73 -331 77 -327
rect 36 -400 40 -396
rect 44 -400 48 -396
rect -41 -483 -37 -479
rect -33 -483 -29 -479
rect -8 -500 0 -489
rect 12 -500 16 -489
rect 24 -502 28 -491
rect 34 -502 42 -493
rect 48 -500 52 -489
rect 60 -502 64 -491
rect 80 -500 88 -489
rect -2 -610 4 -603
rect 33 -608 38 -601
rect 65 -614 69 -610
rect 73 -614 77 -610
rect 36 -672 40 -668
rect 44 -672 48 -668
rect -41 -755 -37 -751
rect -33 -755 -29 -751
rect -8 -772 0 -761
rect 12 -772 16 -761
rect 24 -774 28 -763
rect 34 -774 42 -765
rect 48 -772 52 -761
rect 60 -774 64 -763
rect 80 -772 88 -761
rect -2 -882 4 -875
rect 33 -880 38 -873
rect 65 -886 69 -882
rect 73 -886 77 -882
<< pdcontact >>
rect 36 -99 40 -91
rect 44 -99 48 -91
rect 2 -159 6 -153
rect 34 -162 42 -154
rect 70 -159 74 -153
rect -41 -182 -37 -174
rect -33 -182 -29 -174
rect -2 -279 3 -274
rect 16 -283 22 -277
rect 36 -279 41 -274
rect 65 -313 69 -305
rect 73 -313 77 -305
rect 36 -382 40 -374
rect 44 -382 48 -374
rect 2 -442 6 -436
rect 34 -445 42 -437
rect 70 -442 74 -436
rect -41 -465 -37 -457
rect -33 -465 -29 -457
rect -2 -562 3 -557
rect 16 -566 22 -560
rect 36 -562 41 -557
rect 65 -596 69 -588
rect 73 -596 77 -588
rect 36 -654 40 -646
rect 44 -654 48 -646
rect 2 -714 6 -708
rect 34 -717 42 -709
rect 70 -714 74 -708
rect -41 -737 -37 -729
rect -33 -737 -29 -729
rect -2 -834 3 -829
rect 16 -838 22 -832
rect 36 -834 41 -829
rect 65 -868 69 -860
rect 73 -868 77 -860
<< polysilicon >>
rect 41 -91 43 -88
rect 41 -113 43 -99
rect 41 -120 43 -117
rect 7 -153 11 -148
rect 29 -153 33 -148
rect 43 -153 47 -148
rect 65 -153 69 -148
rect -36 -174 -34 -171
rect 7 -175 11 -162
rect 29 -175 33 -162
rect 9 -179 11 -175
rect 31 -179 33 -175
rect -36 -196 -34 -182
rect -36 -203 -34 -200
rect 7 -206 11 -179
rect 29 -206 33 -179
rect 43 -170 47 -162
rect 65 -170 69 -162
rect 43 -174 45 -170
rect 65 -174 67 -170
rect 43 -206 47 -174
rect 65 -206 69 -174
rect 7 -224 11 -219
rect 29 -224 33 -219
rect 43 -224 47 -219
rect 65 -224 69 -219
rect 7 -274 12 -271
rect 25 -274 30 -271
rect 7 -309 12 -283
rect 7 -318 12 -314
rect 25 -300 30 -283
rect 70 -305 72 -302
rect 25 -318 30 -305
rect 70 -327 72 -313
rect 7 -330 12 -327
rect 25 -330 30 -327
rect 70 -334 72 -331
rect 41 -374 43 -371
rect 41 -396 43 -382
rect 41 -403 43 -400
rect 7 -436 11 -431
rect 29 -436 33 -431
rect 43 -436 47 -431
rect 65 -436 69 -431
rect -36 -457 -34 -454
rect 7 -458 11 -445
rect 29 -458 33 -445
rect 9 -462 11 -458
rect 31 -462 33 -458
rect -36 -479 -34 -465
rect -36 -486 -34 -483
rect 7 -489 11 -462
rect 29 -489 33 -462
rect 43 -453 47 -445
rect 65 -453 69 -445
rect 43 -457 45 -453
rect 65 -457 67 -453
rect 43 -489 47 -457
rect 65 -489 69 -457
rect 7 -507 11 -502
rect 29 -507 33 -502
rect 43 -507 47 -502
rect 65 -507 69 -502
rect 7 -557 12 -554
rect 25 -557 30 -554
rect 7 -592 12 -566
rect 7 -601 12 -597
rect 25 -583 30 -566
rect 70 -588 72 -585
rect 25 -601 30 -588
rect 70 -610 72 -596
rect 7 -613 12 -610
rect 25 -613 30 -610
rect 70 -617 72 -614
rect 41 -646 43 -643
rect 41 -668 43 -654
rect 41 -675 43 -672
rect 7 -708 11 -703
rect 29 -708 33 -703
rect 43 -708 47 -703
rect 65 -708 69 -703
rect -36 -729 -34 -726
rect 7 -730 11 -717
rect 29 -730 33 -717
rect 9 -734 11 -730
rect 31 -734 33 -730
rect -36 -751 -34 -737
rect -36 -758 -34 -755
rect 7 -761 11 -734
rect 29 -761 33 -734
rect 43 -725 47 -717
rect 65 -725 69 -717
rect 43 -729 45 -725
rect 65 -729 67 -725
rect 43 -761 47 -729
rect 65 -761 69 -729
rect 7 -779 11 -774
rect 29 -779 33 -774
rect 43 -779 47 -774
rect 65 -779 69 -774
rect 7 -829 12 -826
rect 25 -829 30 -826
rect 7 -864 12 -838
rect 7 -873 12 -869
rect 25 -855 30 -838
rect 70 -860 72 -857
rect 25 -873 30 -860
rect 70 -882 72 -868
rect 7 -885 12 -882
rect 25 -885 30 -882
rect 70 -889 72 -886
<< polycontact >>
rect 37 -110 41 -106
rect 5 -179 9 -175
rect 27 -179 31 -175
rect -40 -193 -36 -189
rect 45 -174 49 -170
rect 67 -174 71 -170
rect 7 -314 12 -309
rect 25 -305 30 -300
rect 66 -324 70 -320
rect 37 -393 41 -389
rect 5 -462 9 -458
rect 27 -462 31 -458
rect -40 -476 -36 -472
rect 45 -457 49 -453
rect 67 -457 71 -453
rect 7 -597 12 -592
rect 25 -588 30 -583
rect 66 -607 70 -603
rect 37 -665 41 -661
rect 5 -734 9 -730
rect 27 -734 31 -730
rect -40 -748 -36 -744
rect 45 -729 49 -725
rect 67 -729 71 -725
rect 7 -869 12 -864
rect 25 -860 30 -855
rect 66 -879 70 -875
<< metal1 >>
rect 30 -85 88 -81
rect 36 -91 40 -85
rect 44 -106 48 -99
rect 26 -110 37 -106
rect 44 -110 54 -106
rect 44 -113 48 -110
rect 36 -121 40 -117
rect 32 -126 54 -121
rect 83 -130 88 -85
rect -12 -134 88 -130
rect -12 -164 -8 -134
rect 2 -153 6 -134
rect 70 -153 74 -134
rect -47 -168 -8 -164
rect -41 -174 -37 -168
rect -33 -189 -29 -182
rect -15 -179 5 -175
rect 23 -179 27 -175
rect 34 -177 42 -162
rect 49 -174 55 -170
rect 71 -174 75 -170
rect -15 -189 -11 -179
rect 34 -185 96 -177
rect 80 -189 88 -185
rect -51 -193 -40 -189
rect -33 -193 -11 -189
rect -33 -196 -29 -193
rect -8 -197 88 -189
rect -41 -204 -37 -200
rect -54 -208 -28 -204
rect -8 -206 0 -197
rect 12 -203 52 -200
rect 12 -206 16 -203
rect 48 -206 52 -203
rect 24 -227 28 -219
rect -22 -231 28 -227
rect 80 -206 88 -197
rect -22 -247 -17 -231
rect 34 -235 42 -219
rect 60 -227 64 -219
rect 60 -231 110 -227
rect -6 -236 84 -235
rect 0 -241 84 -236
rect -6 -242 84 -241
rect 105 -247 110 -231
rect -22 -251 110 -247
rect -12 -263 59 -258
rect -2 -274 3 -263
rect 36 -274 41 -263
rect 16 -292 22 -283
rect 16 -297 38 -292
rect 18 -305 25 -300
rect 33 -309 38 -297
rect 55 -295 59 -263
rect 55 -299 83 -295
rect 65 -305 69 -299
rect 0 -314 7 -309
rect 33 -314 56 -309
rect 33 -318 38 -314
rect 53 -320 56 -314
rect 73 -320 77 -313
rect 53 -324 66 -320
rect 73 -324 87 -320
rect 73 -327 77 -324
rect -2 -334 4 -327
rect -12 -335 50 -334
rect 65 -335 69 -331
rect -12 -339 83 -335
rect 30 -368 88 -364
rect 36 -374 40 -368
rect 44 -389 48 -382
rect 26 -393 37 -389
rect 44 -393 54 -389
rect 44 -396 48 -393
rect 36 -404 40 -400
rect 32 -409 54 -404
rect 83 -413 88 -368
rect -12 -417 88 -413
rect -12 -447 -8 -417
rect 2 -436 6 -417
rect 70 -436 74 -417
rect -47 -451 -8 -447
rect -41 -457 -37 -451
rect -33 -472 -29 -465
rect -15 -462 5 -458
rect 23 -462 27 -458
rect 34 -460 42 -445
rect 49 -457 55 -453
rect 71 -457 75 -453
rect -15 -472 -11 -462
rect 34 -468 96 -460
rect 80 -472 88 -468
rect -51 -476 -40 -472
rect -33 -476 -11 -472
rect -33 -479 -29 -476
rect -8 -480 88 -472
rect -41 -487 -37 -483
rect -54 -491 -28 -487
rect -8 -489 0 -480
rect 12 -486 52 -483
rect 12 -489 16 -486
rect 48 -489 52 -486
rect 24 -510 28 -502
rect -22 -514 28 -510
rect 80 -489 88 -480
rect -22 -530 -17 -514
rect 34 -518 42 -502
rect 60 -510 64 -502
rect 60 -514 110 -510
rect -6 -519 84 -518
rect 0 -524 84 -519
rect -6 -525 84 -524
rect 105 -530 110 -514
rect -22 -534 110 -530
rect -12 -546 59 -541
rect -2 -557 3 -546
rect 36 -557 41 -546
rect 16 -575 22 -566
rect 16 -580 38 -575
rect 18 -588 25 -583
rect 33 -592 38 -580
rect 55 -578 59 -546
rect 55 -582 83 -578
rect 65 -588 69 -582
rect 0 -597 7 -592
rect 33 -597 56 -592
rect 33 -601 38 -597
rect 53 -603 56 -597
rect 73 -603 77 -596
rect 53 -607 66 -603
rect 73 -607 87 -603
rect 73 -610 77 -607
rect -2 -617 4 -610
rect -12 -618 50 -617
rect 65 -618 69 -614
rect -12 -622 83 -618
rect 30 -640 88 -636
rect 36 -646 40 -640
rect 44 -661 48 -654
rect 26 -665 37 -661
rect 44 -665 54 -661
rect 44 -668 48 -665
rect 36 -676 40 -672
rect 32 -681 54 -676
rect 83 -685 88 -640
rect -12 -689 88 -685
rect -12 -719 -8 -689
rect 2 -708 6 -689
rect 70 -708 74 -689
rect -47 -723 -8 -719
rect -41 -729 -37 -723
rect -33 -744 -29 -737
rect -15 -734 5 -730
rect 23 -734 27 -730
rect 34 -732 42 -717
rect 49 -729 55 -725
rect 71 -729 75 -725
rect -15 -744 -11 -734
rect 34 -740 96 -732
rect 80 -744 88 -740
rect -51 -748 -40 -744
rect -33 -748 -11 -744
rect -33 -751 -29 -748
rect -8 -752 88 -744
rect -41 -759 -37 -755
rect -54 -763 -28 -759
rect -8 -761 0 -752
rect 12 -758 52 -755
rect 12 -761 16 -758
rect 48 -761 52 -758
rect 24 -782 28 -774
rect -22 -786 28 -782
rect 80 -761 88 -752
rect -22 -802 -17 -786
rect 34 -790 42 -774
rect 60 -782 64 -774
rect 60 -786 110 -782
rect -6 -791 84 -790
rect 0 -796 84 -791
rect -6 -797 84 -796
rect 105 -802 110 -786
rect -22 -806 110 -802
rect -12 -818 59 -813
rect -2 -829 3 -818
rect 36 -829 41 -818
rect 16 -847 22 -838
rect 16 -852 38 -847
rect 18 -860 25 -855
rect 33 -864 38 -852
rect 55 -850 59 -818
rect 55 -854 83 -850
rect 65 -860 69 -854
rect 0 -869 7 -864
rect 33 -869 56 -864
rect 33 -873 38 -869
rect 53 -875 56 -869
rect 73 -875 77 -868
rect 53 -879 66 -875
rect 73 -879 87 -875
rect 73 -882 77 -879
rect -2 -889 4 -882
rect -12 -890 50 -889
rect 65 -890 69 -886
rect -12 -894 83 -890
<< m2contact >>
rect 54 -110 60 -105
rect 55 -174 60 -169
rect -59 -208 -54 -203
rect -28 -208 -23 -203
rect -6 -241 0 -236
rect 54 -393 60 -388
rect 55 -457 60 -452
rect -59 -491 -54 -486
rect -28 -491 -23 -486
rect -6 -524 0 -519
rect 54 -665 60 -660
rect 55 -729 60 -724
rect -59 -763 -54 -758
rect -28 -763 -23 -758
rect -6 -796 0 -791
<< metal2 >>
rect -59 -203 -54 -126
rect 55 -169 60 -110
rect -28 -236 -23 -208
rect -28 -241 -6 -236
rect -59 -486 -54 -409
rect 55 -452 60 -393
rect -28 -519 -23 -491
rect -28 -524 -6 -519
rect -59 -758 -54 -681
rect 55 -724 60 -665
rect -28 -791 -23 -763
rect -28 -796 -6 -791
<< m3contact >>
rect -59 -126 -54 -121
rect -59 -409 -54 -404
rect -59 -681 -54 -676
<< m123contact >>
rect 27 -126 32 -121
rect 27 -409 32 -404
rect 27 -681 32 -676
<< metal3 >>
rect -54 -126 27 -121
rect -54 -409 27 -404
rect -54 -681 27 -676
use XORinv  XORinv_0
timestamp 1638834489
transform 1 0 -22 0 1 28
box -37 0 132 170
use AND2  AND2_0
timestamp 1638834295
transform 1 0 13 0 1 0
box -25 -60 74 21
<< labels >>
rlabel metal1 -47 -208 -23 -204 1 gnd
rlabel metal1 37 -239 37 -239 1 gnd
rlabel metal1 38 -132 38 -132 5 vdd
rlabel metal1 59 -582 83 -578 5 vdd
rlabel metal1 38 -415 38 -415 5 vdd
rlabel metal1 37 -522 37 -522 1 gnd
rlabel metal1 -47 -491 -23 -487 1 gnd
rlabel metal1 -47 -451 -23 -447 5 vdd
rlabel metal1 59 -854 83 -850 5 vdd
rlabel metal1 38 -687 38 -687 5 vdd
rlabel metal1 37 -794 37 -794 1 gnd
rlabel metal1 -47 -763 -23 -759 1 gnd
rlabel metal1 -47 -723 -23 -719 5 vdd
rlabel metal1 30 -640 54 -636 5 vdd
rlabel metal1 27 -126 54 -121 1 gnd
rlabel metal1 27 -409 54 -404 1 gnd
rlabel polycontact 5 -179 9 -175 1 b2bar
rlabel polycontact 27 -179 31 -175 1 a2
rlabel polycontact 45 -174 49 -170 1 a2bar
rlabel polycontact 67 -174 71 -170 1 b2
rlabel metal1 0 -314 12 -309 1 a2
rlabel metal1 88 -185 96 -177 1 p2
rlabel metal1 83 -324 87 -320 1 g2
rlabel space 0 -35 12 -30 1 a3
rlabel metal1 0 -597 12 -592 1 a1
rlabel polycontact 5 -462 9 -458 1 b1bar
rlabel polycontact 27 -462 31 -458 1 a1
rlabel polycontact 45 -457 49 -453 1 a1bar
rlabel polycontact 67 -457 71 -453 1 b1
rlabel metal1 88 -468 96 -460 1 p1
rlabel metal1 83 -607 87 -603 1 g1
rlabel metal1 88 -740 96 -732 1 p0
rlabel metal1 83 -879 87 -875 1 g0
rlabel metal1 0 -869 12 -864 1 a0
rlabel polycontact 5 -734 9 -730 1 b0bar
rlabel polycontact -40 -748 -36 -744 1 b0
rlabel polycontact 67 -729 71 -725 1 b0
rlabel polycontact 45 -729 49 -725 1 a0bar
rlabel polycontact 27 -734 31 -730 1 a0
rlabel metal1 38 -892 38 -892 1 gnd
rlabel polycontact 37 -665 41 -661 1 a0
rlabel m2contact 54 -665 60 -660 1 a0bar
rlabel metal1 33 -620 33 -620 1 gnd
rlabel metal1 23 -544 23 -544 1 vdd
rlabel polycontact -40 -476 -36 -472 1 b1
rlabel polycontact 37 -393 41 -389 1 a1
rlabel metal1 47 -366 47 -366 1 vdd
rlabel metal1 32 -337 32 -337 1 gnd
rlabel metal1 44 -261 44 -261 1 vdd
rlabel polycontact -40 -193 -36 -189 1 b2
rlabel polycontact 37 -110 41 -106 1 a2
rlabel space 5 100 9 104 1 b3bar
rlabel space 27 100 31 104 1 a3
rlabel space 45 105 49 109 1 a3bar
rlabel space 67 105 71 109 1 b3
rlabel space 88 94 96 102 1 p3
rlabel space 83 -45 87 -41 1 g3
rlabel polycontact 66 -324 70 -320 1 g2in
rlabel polycontact 66 -607 70 -603 1 g1in
rlabel polycontact 66 -879 70 -875 1 g0in
rlabel space 66 -45 70 -41 1 g3in
rlabel space 18 -27 30 -22 1 b3
rlabel metal1 18 -305 30 -300 1 b2
rlabel metal1 18 -588 30 -583 1 b1
rlabel metal1 20 -816 20 -816 1 vdd
rlabel metal1 18 -860 30 -855 1 b0
<< end >>
