* Full Adder pre-simulation

.include TSMC_180nm.txt
.include NOT_SUB.sub
.include AND2.sub
.include AND3.sub
.include AND4.sub
.include AND5.sub
.include XOR.sub
.include OR.sub

.param LAMBDA = 0.18u
.param width_N = {10*LAMBDA}
.param width_P = {2.5*width_N}

vdd vdd gnd 2.0V

Vin1 A gnd pulse(0 2.0 0 0.01p 0.01p 10n 20n)
Vin2 B gnd pulse(0 2.0 0 0.01p 0.01p 20n 40n)
Vin3 C gnd pulse(0 2.0 0 0.01p 0.01p 40n 80n)


xG1 A B P XOR
xG2 A B G AND2

xG3 C P sum XOR
xG4 P C Cx AND2

xG5 Cx G Cplus OR

.control
tran 1n 120n
plot v(A)
plot v(B)
plot v(C)
plot v(sum)
plot v(Cplus)
.endc
.end