* SPICE3 file created from AND3.ext - technology: scmos

.include TSMC_180nm.txt

vdd vdd gnd 2.0V

.option scale=0.09u

Vin1 A gnd pulse(0 2.0 0 0.01p 0.01p 10n 20n)
Vin2 B gnd pulse(0 2.0 0 0.01p 0.01p 20n 40n)
Vin3 C gnd pulse(0 2.0 0 0.01p 0.01p 40n 80n)

M1000 outout OUT vdd NOT_0/w_0_0# CMOSP w=8 l=2
+  ad=40 pd=26 as=112 ps=74
M1001 outout OUT gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=42 ps=38
M1002 OUT A vdd w_n32_7# CMOSP w=6 l=2
+  ad=78 pd=50 as=0 ps=0
M1003 vdd B OUT w_n32_7# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_n10_n22# B a_n18_n22# gnd CMOSN w=3 l=2
+  ad=18 pd=18 as=18 ps=18
M1005 OUT A a_n10_n22# gnd CMOSN w=3 l=2
+  ad=25 pd=22 as=0 ps=0
M1006 a_n18_n22# C gnd gnd CMOSN w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 OUT C vdd w_n32_7# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0

.control
tran 1n 160n
plot v(A) 
plot v(B)
plot v(C)
plot v(outout)
.endc
.end