magic
tech scmos
timestamp 1638851182
<< metal1 >>
rect 285 917 612 918
rect 285 908 776 917
rect 285 853 290 908
rect 447 907 776 908
rect 142 849 290 853
rect 170 754 236 759
rect 489 738 711 742
rect 173 626 201 631
rect 206 626 235 631
rect 184 618 216 623
rect 752 591 776 907
rect 723 587 955 591
rect 142 570 150 574
rect 146 542 150 570
rect 184 553 205 556
rect 184 552 200 553
rect 146 537 173 542
rect 167 510 173 537
rect 167 503 585 510
rect 190 447 197 503
rect 752 463 776 587
rect 752 456 802 463
rect 208 438 214 440
rect 208 436 210 438
rect 207 431 210 432
rect 184 428 210 431
rect 184 427 208 428
rect 210 416 214 417
rect 190 369 197 408
rect 179 362 197 369
rect 168 291 173 327
rect 142 287 173 291
rect 179 267 186 362
rect 810 361 811 369
rect 198 344 201 348
rect 206 348 210 349
rect 206 345 211 348
rect 198 302 203 344
rect 918 337 961 341
rect 198 298 208 302
rect 203 259 208 298
rect 203 254 222 259
<< m2contact >>
rect 147 988 155 996
rect 382 802 390 810
rect 711 737 723 742
rect 147 709 155 717
rect 168 626 173 631
rect 201 626 206 631
rect 177 618 184 623
rect 585 610 593 618
rect 711 587 723 592
rect 177 552 184 557
rect 693 546 698 551
rect 585 502 593 510
rect 802 456 810 463
rect 190 441 197 447
rect 203 436 208 441
rect 177 427 184 432
rect 190 408 197 413
rect 168 327 173 332
rect 802 361 810 369
rect 201 344 206 349
rect 210 337 215 342
rect 912 337 918 342
rect 208 328 213 333
rect 179 262 186 267
rect 238 262 243 267
<< metal2 >>
rect 155 988 194 996
rect 155 709 184 717
rect 176 635 184 709
rect 168 332 173 626
rect 177 623 184 635
rect 177 557 184 618
rect 177 432 184 552
rect 188 519 194 988
rect 382 701 390 802
rect 201 696 390 701
rect 201 631 206 696
rect 188 512 208 519
rect 177 340 184 427
rect 190 413 197 441
rect 203 441 208 512
rect 585 510 593 610
rect 711 592 722 737
rect 698 546 918 550
rect 203 434 208 436
rect 203 349 207 434
rect 802 369 810 456
rect 912 342 918 546
rect 177 337 210 340
rect 177 336 203 337
rect 173 328 208 332
rect 186 262 238 267
<< m123contact >>
rect 165 754 170 759
rect 149 427 155 433
rect 203 545 208 550
rect 211 420 216 425
<< metal3 >>
rect 165 611 170 754
rect 157 607 170 611
rect 157 549 163 607
rect 157 545 203 549
rect 157 433 163 545
rect 155 427 163 433
rect 157 424 163 427
rect 157 420 211 424
use PandG  PandG_0
timestamp 1638851043
transform 1 0 59 0 1 894
box -59 -894 110 198
use XORinv  XORinv_3
timestamp 1638850046
transform 1 0 982 0 1 945
box -37 0 132 170
use CLA  CLA_0
timestamp 1638851043
transform 1 0 238 0 1 725
box -35 -496 679 152
use XORinv  XORinv_0
timestamp 1638850046
transform 1 0 984 0 1 725
box -37 0 132 170
use XORinv  XORinv_1
timestamp 1638850046
transform 1 0 984 0 1 529
box -37 0 132 170
use XORinv  XORinv_2
timestamp 1638850046
transform 1 0 988 0 1 279
box -37 0 132 170
<< labels >>
rlabel space 1015 351 1019 355 1 c3bar
rlabel space 1037 351 1041 355 1 p3
rlabel space 1047 420 1051 424 1 p3
rlabel space 1055 356 1059 360 1 p3bar
rlabel space 1077 356 1081 360 1 c3
rlabel space 1011 601 1015 605 1 c2bar
rlabel space 1033 601 1037 605 1 p2
rlabel space 1051 606 1055 610 1 p2bar
rlabel space 1043 670 1047 674 1 p2
rlabel space 1073 606 1077 610 1 c2
rlabel space 966 783 970 787 1 c1
rlabel space 1073 802 1077 806 1 c1
rlabel space 1011 797 1015 801 1 c1bar
rlabel space 1033 797 1037 801 1 p1
rlabel space 1051 802 1055 806 1 p1bar
rlabel space 1043 866 1047 870 1 p1
rlabel space 964 1003 968 1007 1 c0
rlabel space 1009 1017 1013 1021 1 c0bar
rlabel space 1031 1017 1035 1021 1 p0
rlabel space 1049 1022 1053 1026 1 p0bar
rlabel space 1041 1086 1045 1090 1 p0
rlabel space 1071 1022 1075 1026 1 c0
<< end >>
