* Carry-lookahead adder for 4 bit inputs

.include TSMC_180nm.txt
.include NOT_SUB.sub
.include AND2.sub
.include AND3.sub
.include AND4.sub
.include AND5.sub
.include XOR.sub
.include OR.sub
.include PROP_GEN.sub
.include CLA.sub
.include SUMMER.sub

.param LAMBDA = 0.18u
.param width_N = {10*LAMBDA}
.param width_P = {2.5*width_N}

* Defining the inputs
vdd vdd gnd 2.0V

Vin1 A0 gnd pulse(2.0 0 0ns 100ps 100ps 10ns 20ns)
Vin2 A1 gnd pulse(0 2.0 0ns 100ps 100ps 20ns 40ns)
Vin3 A2 gnd pulse(0 2.0 0ns 100ps 100ps 20ns 40ns)
Vin4 A3 gnd pulse(0 2.0 0ns 100ps 100ps 20ns 40ns)

Vin5 B0 gnd pulse(2.0 0 0ns 100ps 100ps 20ns 40ns)
Vin6 B1 gnd pulse(0 2.0 0ns 100ps 100ps 20ns 40ns)
Vin7 B2 gnd pulse(0 2.0 0ns 100ps 100ps 20ns 40ns)
Vin8 B3 gnd pulse(0 2.0 0ns 100ps 100ps 20ns 40ns)

Vin9 C0 gnd pulse(0 2.0 0ns 100ps 100ps 40ns 80ns)

* Making the logic part

* Generating the propogate and generate of the carry-lookahead adder
xG1 A0 B0 A1 B1 A2 B2 A3 B3 P0 G0 P1 G1 P2 G2 P3 G3 PROP_GEN

* Generating the carry bits of the carry-lookahead adder
xG2 C0 P0 G0 G1 P1 G2 P2 G3 P3 C1 C2 C3 C4 CLA

* Generating the sums of the carry-lookahead adder
xG3 P0 P1 P2 P3 C0 C1 C2 C3 S0 S1 S2 S3 SUMMER

* Plotting the inputs and outputs
.control
tran 1n 80n
set curplottitle= Aditya-Nair-2020102022-3-Final
plot v(S0)
plot v(S1)
plot v(S2)
plot v(S3)
plot v(C4)
.endc
.end