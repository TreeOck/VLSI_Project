magic
tech scmos
timestamp 1638828285
<< nwell >>
rect -25 -47 83 1
<< ntransistor >>
rect -7 -113 0 -92
rect 53 -113 60 -92
<< ptransistor >>
rect -7 -35 0 -9
rect 53 -35 60 -9
<< ndiffusion >>
rect -25 -102 -7 -92
rect -25 -108 -21 -102
rect -13 -108 -7 -102
rect -25 -113 -7 -108
rect 0 -100 53 -92
rect 0 -106 20 -100
rect 30 -106 53 -100
rect 0 -113 53 -106
rect 60 -102 83 -92
rect 60 -108 68 -102
rect 76 -108 83 -102
rect 60 -113 83 -108
<< pdiffusion >>
rect -18 -18 -7 -9
rect -18 -24 -17 -18
rect -9 -24 -7 -18
rect -18 -35 -7 -24
rect 0 -35 53 -9
rect 60 -20 75 -9
rect 60 -26 64 -20
rect 72 -26 75 -20
rect 60 -35 75 -26
<< ndcontact >>
rect -21 -108 -13 -102
rect 20 -106 30 -100
rect 68 -108 76 -102
<< pdcontact >>
rect -17 -24 -9 -18
rect 64 -26 72 -20
<< polysilicon >>
rect -7 -9 0 6
rect 53 -9 60 6
rect -7 -50 0 -35
rect -7 -92 0 -58
rect 53 -50 60 -35
rect 53 -92 60 -58
rect -7 -117 0 -113
rect 53 -117 60 -113
rect 127 -122 131 -118
<< polycontact >>
rect -7 -58 0 -50
rect 53 -58 60 -50
<< metal1 >>
rect -24 12 118 17
rect -17 -18 -9 12
rect -18 -58 -7 -50
rect 42 -58 53 -50
rect 64 -65 72 -26
rect 20 -73 97 -65
rect 20 -100 30 -73
rect -21 -133 -13 -108
rect 68 -133 76 -108
rect 92 -118 97 -73
rect 113 -93 118 12
rect 113 -97 122 -93
rect 92 -122 116 -118
rect -21 -137 122 -133
rect -21 -139 144 -137
use NOTNOT  NOTNOT_0
timestamp 1638796604
transform 1 0 120 0 1 -117
box -4 -20 28 24
<< end >>
