magic
tech scmos
timestamp 1638843228
<< nwell >>
rect -32 7 11 25
<< ntransistor >>
rect -20 -22 -18 -19
rect -12 -22 -10 -19
rect -4 -22 -2 -19
<< ptransistor >>
rect -20 13 -18 19
rect -12 13 -10 19
rect -4 13 -2 19
<< ndiffusion >>
rect -22 -22 -20 -19
rect -18 -22 -12 -19
rect -10 -22 -4 -19
rect -2 -22 1 -19
<< pdiffusion >>
rect -22 13 -20 19
rect -18 13 -17 19
rect -13 13 -12 19
rect -10 13 -9 19
rect -5 13 -4 19
rect -2 13 1 19
<< ndcontact >>
rect -26 -23 -22 -19
rect 1 -22 5 -18
<< pdcontact >>
rect -26 13 -22 19
rect -17 13 -13 19
rect -9 13 -5 19
rect 1 13 5 19
<< polysilicon >>
rect -20 19 -18 22
rect -12 19 -10 22
rect -4 19 -2 22
rect -20 -12 -18 13
rect -12 -5 -10 13
rect -4 3 -2 13
rect -20 -19 -18 -16
rect -12 -19 -10 -9
rect -4 -19 -2 -1
rect -20 -25 -18 -22
rect -12 -25 -10 -22
rect -4 -25 -2 -22
<< polycontact >>
rect -6 -1 -2 3
rect -14 -9 -10 -5
rect -22 -16 -18 -12
<< metal1 >>
rect -32 28 21 32
rect -26 19 -22 28
rect -9 19 -5 28
rect -17 9 -13 13
rect 1 9 5 13
rect 17 10 21 28
rect -17 6 5 9
rect -32 -1 -6 3
rect 1 -2 5 6
rect -32 -9 -14 -5
rect 1 -6 17 -2
rect -32 -16 -22 -12
rect 1 -18 5 -6
rect 13 -15 17 -6
rect -26 -26 -22 -23
rect -32 -30 21 -26
use NOT  NOT_0
timestamp 1638826985
transform 1 0 21 0 1 -10
box -4 -20 28 24
<< labels >>
rlabel metal1 -12 -30 -7 -26 1 gnd
rlabel metal1 9 -4 9 -4 1 out1
rlabel metal1 -6 30 -6 30 5 vdd
<< end >>
