* NOT gate pre-simulation

.include TSMC_180nm.txt

.param LAMBDA = 0.18u
.param width_N = {10*LAMBDA}
.param width_P = {2.5*width_N}

vdd vdd gnd 2.0V

Vin A gnd pulse(0 2.0 0 0.01p 0.01p 10n 20n)

M1 B A vdd vdd CMOSP W={width_P} L={LAMBDA}
+ AS = {5*width_P*LAMBDA} PS = {10*LAMBDA + 2*width_P} AD = {5*width_P*LAMBDA} PD = {10*LAMBDA + 2*width_P}

M2 B A gnd gnd CMOSN W={width_N} L={LAMBDA}
+ AS = {5*width_N*LAMBDA} PS = {10*LAMBDA + 2*width_N} AD = {5*width_N*LAMBDA} PD = {10*LAMBDA + 2*width_N}

.control
tran 1n 100n
set curplottitle= Aditya-Nair-2020102022-3-NOT
plot v(A) 
plot v(B)
.endc
.end
