* AND gate pre-simulation

.include TSMC_180nm.txt
.include NOT_SUB.sub

.param LAMBDA = 0.18u
.param width_N = {10*LAMBDA}
.param width_P = {2.5*width_N}

vdd Vcc GND 2.0V

Vin1 A GND pulse(0 2.0 0 0.01p 0.01p 10n 20n)
Vin2 B GND pulse(0 2.0 0 0.01p 0.01p 20n 40n)

M1 C A Vcc Vcc CMOSP W={width_P} L={LAMBDA}
+ AS = {5*width_P*LAMBDA} PS = {10*LAMBDA + 2*width_P} AD = {5*width_P*LAMBDA} PD = {10*LAMBDA + 2*width_P}

M2 C B Vcc Vcc CMOSP W={width_P} L={LAMBDA}
+ AS = {5*width_P*LAMBDA} PS = {10*LAMBDA + 2*width_P} AD = {5*width_P*LAMBDA} PD = {10*LAMBDA + 2*width_P}

M3 C B D D CMOSN W={width_N} L={LAMBDA}
+ AS = {5*width_N*LAMBDA} PS = {10*LAMBDA + 2*width_N} AD = {5*width_N*LAMBDA} PD = {10*LAMBDA + 2*width_N}

M4 D A GND GND CMOSN W={width_N} L={LAMBDA}
+ AS = {5*width_N*LAMBDA} PS = {10*LAMBDA + 2*width_N} AD = {5*width_N*LAMBDA} PD = {10*LAMBDA + 2*width_N}

xG1 C E NOTNOT

.control
tran 1n 120n
set curplottitle= Aditya-Nair-2020102022-3-AND2
plot v(A) 
plot v(B)
plot v(C)
plot v(E)
.endc

.end