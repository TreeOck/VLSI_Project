magic
tech scmos
timestamp 1638844744
<< nwell >>
rect -6 -6 46 12
<< ntransistor >>
rect 5 -52 7 -46
rect 15 -52 17 -46
rect 23 -52 25 -46
rect 32 -52 34 -46
<< ptransistor >>
rect 5 0 7 6
rect 15 0 17 6
rect 23 0 25 6
rect 32 0 34 6
<< ndiffusion >>
rect 4 -52 5 -46
rect 7 -52 15 -46
rect 17 -52 23 -46
rect 25 -52 32 -46
rect 34 -52 37 -46
<< pdiffusion >>
rect 4 0 5 6
rect 7 0 9 6
rect 13 0 15 6
rect 17 0 18 6
rect 22 0 23 6
rect 25 0 27 6
rect 31 0 32 6
rect 34 0 35 6
rect 39 0 40 6
<< ndcontact >>
rect 0 -52 4 -46
rect 37 -52 41 -46
<< pdcontact >>
rect 0 0 4 6
rect 9 0 13 6
rect 18 0 22 6
rect 27 0 31 6
rect 35 0 39 6
<< polysilicon >>
rect 5 6 7 9
rect 15 6 17 9
rect 23 6 25 9
rect 32 6 34 9
rect 5 -16 7 0
rect 5 -46 7 -20
rect 15 -25 17 0
rect 15 -46 17 -29
rect 23 -32 25 0
rect 23 -46 25 -36
rect 32 -39 34 0
rect 32 -46 34 -43
rect 5 -55 7 -52
rect 15 -55 17 -52
rect 23 -55 25 -52
rect 32 -55 34 -52
<< polycontact >>
rect 3 -20 7 -16
rect 13 -29 17 -25
rect 21 -36 25 -32
rect 30 -43 34 -39
<< metal1 >>
rect -6 18 53 22
rect 0 6 4 18
rect 18 6 22 18
rect 35 6 39 18
rect 9 -11 13 0
rect 27 -11 31 0
rect 9 -13 41 -11
rect 10 -15 41 -13
rect -6 -20 3 -16
rect -6 -24 3 -23
rect -6 -25 6 -24
rect -6 -27 13 -25
rect 3 -29 13 -27
rect 37 -31 41 -15
rect 49 -28 53 18
rect -6 -36 21 -32
rect 37 -35 49 -31
rect -6 -43 30 -39
rect 37 -46 41 -35
rect 0 -64 4 -52
rect 45 -53 49 -35
rect -6 -68 53 -64
use NOT  NOT_0
timestamp 1638826985
transform 1 0 53 0 1 -48
box -4 -20 28 24
<< labels >>
rlabel metal1 22 20 22 20 5 vdd
rlabel metal1 42 -33 42 -33 1 out1
rlabel metal1 20 -66 20 -66 1 gnd
<< end >>
