* SPICE3 file created from AND4.ext - technology: scmos

.include TSMC_180nm.txt

vdd vdd gnd 2.0V

.option scale=0.09u

Vin1 A gnd pulse(0 2.0 0 0.01p 0.01p 10n 20n)
Vin2 B gnd pulse(0 2.0 0 0.01p 0.01p 20n 40n)
Vin3 C gnd pulse(0 2.0 0 0.01p 0.01p 40n 80n)
Vin4 D gnd pulse(0 2.0 0 0.01p 0.01p 80n 160n)

M1000 outout OUT vdd NOT_0/w_0_0# CMOSP w=8 l=2
+  ad=40 pd=26 as=142 ps=96
M1001 outout OUT gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=50 ps=40
M1002 a_7_n52# A gnd gnd CMOSN w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1003 a_25_n52# C a_17_n52# gnd CMOSN w=6 l=2
+  ad=42 pd=26 as=36 ps=24
M1004 vdd B OUT w_n6_n6# CMOSP w=6 l=2
+  ad=0 pd=0 as=90 ps=54
M1005 vdd D OUT w_n6_n6# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 OUT C vdd w_n6_n6# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 OUT D a_25_n52# gnd CMOSN w=6 l=2
+  ad=42 pd=26 as=0 ps=0
M1008 OUT A vdd w_n6_n6# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_17_n52# B a_7_n52# gnd CMOSN w=6 l=2
+  ad=0 pd=0 as=0 ps=0

.control
tran 1n 320n
plot v(A) 
plot v(B)
plot v(C)
plot v(D)
plot v(outout)
.endc
.end