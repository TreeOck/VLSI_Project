magic
tech scmos
timestamp 1638850046
<< metal1 >>
rect 76 166 110 170
rect 75 141 77 145
rect 105 121 110 166
rect 10 117 22 121
rect 102 117 110 121
rect 10 87 14 117
rect -2 83 14 87
rect 71 77 77 81
rect 7 72 23 76
rect 45 72 46 76
rect 7 62 11 72
rect 3 58 11 62
rect -32 43 -24 47
<< m2contact >>
rect 77 141 82 146
rect 77 77 82 82
rect -37 43 -32 48
rect -6 43 -1 48
rect 16 10 22 15
<< metal2 >>
rect -37 48 -32 125
rect 77 82 82 141
rect -6 15 -1 43
rect -6 10 16 15
<< m3contact >>
rect -37 125 -32 130
<< m123contact >>
rect 49 125 54 130
<< metal3 >>
rect -32 125 49 130
use NOT  NOT_1
timestamp 1638826985
transform 1 0 52 0 1 146
box -4 -20 28 24
use NOT  NOT_0
timestamp 1638826985
transform 1 0 -25 0 1 63
box -4 -20 28 24
use XOR  XOR_0
timestamp 1638801340
transform 1 0 74 0 1 86
box -74 -86 58 35
<< end >>
