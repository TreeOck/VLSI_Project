* Combinational circuit-1 pre-simulation

.include TSMC_180nm.txt
.include NOT_SUB.sub
.include AND2.sub
.include AND3.sub
.include AND4.sub
.include AND5.sub
.include XOR.sub
.include OR.sub

.param LAMBDA = 0.18u
.param width_N = {10*LAMBDA}
.param width_P = {2.5*width_N}

vdd vdd gnd 2.0V

Vin1 A0 gnd pulse(0 2.0 0 0.01p 0.01p 10n 20n)
Vin2 B0 gnd pulse(0 2.0 0 0.01p 0.01p 20n 40n)
Vin3 Cin gnd pulse(0 2.0 0 0.01p 0.01p 40n 80n)

xG1 A0 B0 P0 XOR
xG2 A0 B0 G0 AND2

xG3 P0 Cin x1 AND2

xG4 G0 x1 C1 OR

.control
tran 1n 120n
plot v(A0)
plot v(B0)
plot v(Cin)
plot v(P0)
plot v(G0)
plot v(C1)
.endc
.end