magic
tech scmos
timestamp 1638801340
<< nwell >>
rect -57 -3 29 18
<< ntransistor >>
rect -45 -54 -41 -41
rect -23 -54 -19 -41
rect -9 -54 -5 -41
rect 13 -54 17 -41
<< ptransistor >>
rect -45 3 -41 12
rect -23 3 -19 12
rect -9 3 -5 12
rect 13 3 17 12
<< ndiffusion >>
rect -67 -52 -60 -41
rect -52 -52 -45 -41
rect -67 -54 -45 -52
rect -41 -52 -40 -41
rect -36 -43 -23 -41
rect -36 -52 -28 -43
rect -41 -54 -28 -52
rect -24 -54 -23 -43
rect -19 -45 -9 -41
rect -19 -54 -18 -45
rect -10 -54 -9 -45
rect -5 -52 -4 -41
rect 0 -43 13 -41
rect 0 -52 8 -43
rect -5 -54 8 -52
rect 12 -54 13 -43
rect 17 -52 28 -41
rect 36 -52 43 -41
rect 17 -54 43 -52
<< pdiffusion >>
rect -51 6 -50 12
rect -46 6 -45 12
rect -51 3 -45 6
rect -41 3 -23 12
rect -19 11 -9 12
rect -19 3 -18 11
rect -10 3 -9 11
rect -5 3 13 12
rect 17 6 18 12
rect 22 6 23 12
rect 17 3 23 6
<< ndcontact >>
rect -60 -52 -52 -41
rect -40 -52 -36 -41
rect -28 -54 -24 -43
rect -18 -54 -10 -45
rect -4 -52 0 -41
rect 8 -54 12 -43
rect 28 -52 36 -41
<< pdcontact >>
rect -50 6 -46 12
rect -18 3 -10 11
rect 18 6 22 12
<< polysilicon >>
rect -45 12 -41 17
rect -23 12 -19 17
rect -9 12 -5 17
rect 13 12 17 17
rect -45 -10 -41 3
rect -23 -10 -19 3
rect -43 -14 -41 -10
rect -21 -14 -19 -10
rect -45 -41 -41 -14
rect -23 -41 -19 -14
rect -9 -5 -5 3
rect 13 -5 17 3
rect -9 -9 -7 -5
rect 13 -9 15 -5
rect -9 -41 -5 -9
rect 13 -41 17 -9
rect -45 -59 -41 -54
rect -23 -59 -19 -54
rect -9 -59 -5 -54
rect 13 -59 17 -54
<< polycontact >>
rect -47 -14 -43 -10
rect -25 -14 -21 -10
rect -7 -9 -3 -5
rect 15 -9 19 -5
<< metal1 >>
rect -57 31 29 35
rect -50 12 -46 31
rect 18 12 22 31
rect -51 -14 -47 -10
rect -29 -14 -25 -10
rect -18 -12 -10 3
rect -3 -9 1 -5
rect 19 -9 23 -5
rect -18 -20 44 -12
rect 28 -24 36 -20
rect -60 -32 36 -24
rect -60 -41 -52 -32
rect -40 -38 0 -35
rect -40 -41 -36 -38
rect -4 -41 0 -38
rect -28 -62 -24 -54
rect -74 -66 -24 -62
rect 28 -41 36 -32
rect -74 -82 -69 -66
rect -18 -70 -10 -54
rect 8 -62 12 -54
rect 8 -66 58 -62
rect -58 -77 32 -70
rect 53 -82 58 -66
rect -74 -86 58 -82
<< labels >>
rlabel metal1 36 -20 44 -12 1 out
rlabel metal1 -15 -74 -15 -74 1 gnd
rlabel metal1 -14 33 -14 33 5 vdd
<< end >>
